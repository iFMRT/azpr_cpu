﻿/*
 -- ============================================================================
 -- FILE NAME	: uart.v
 -- DESCRIPTION : Universal Asynchronous Receiver and Transmitter
 -- ----------------------------------------------------------------------------
 -- Revision  Date		  Coding_by	 Comment
 -- 1.0.0	  2011/06/27  suito		 ???????
 -- ============================================================================
*/

/********** ?????a???????? **********/
`include "nettype.h"
`include "stddef.h"
`include "global_config.h"

/********** ???e??a???????? **********/
`include "uart.h"

/********** ????`?? **********/
module uart (
	/********** ????a? & ???a? **********/
	input  wire				   clk,		 // ????a?
	input  wire				   reset,	 // ???????a?
	/********** ?刅?????????`?? **********/
	input  wire				   cs_,		 // ???a??????
	input  wire				   as_,		 // ??????????`??
	input  wire				   rw,		 // Read / Write
	input  wire [`UartAddrBus] addr,	 // ?????
	input  wire [`WordDataBus] wr_data,	 // ?????z???`??
	output wire [`WordDataBus] rd_data,	 // ?i???????`??
	output wire				   rdy_,	 // ????
	/********** ????z?? **********/
	output wire				   irq_rx,	 // ???????????z??
	output wire				   irq_tx,	 // ???????????z??
	/********** UART?????????	**********/
	input  wire				   rx,		 // UART???????
	output wire				   tx		 // UART???????
);

	/********** ??????? **********/
	// ????????
	wire					   rx_busy;	 // ?????刅??
	wire					   rx_end;	 // ???????????
	wire [`ByteDataBus]		   rx_data;	 // ?????`??
	// ????????
	wire					   tx_busy;	 // ?????刅??
	wire					   tx_end;	 // ???????????
	wire					   tx_start; // ?????_????
	wire [`ByteDataBus]		   tx_data;	 // ?????`??

	/********** UART????????`?? **********/
	uart_ctrl uart_ctrl (
		/********** ????a? & ???a? **********/
		.clk	  (clk),	   // ????a?
		.reset	  (reset),	   // ???????a?
		/********** Host Interface **********/
		.cs_	  (cs_),	   // ???a??????
		.as_	  (as_),	   // ??????????`??
		.rw		  (rw),		   // Read / Write
		.addr	  (addr),	   // ?????
		.wr_data  (wr_data),   // ?????z???`??
		.rd_data  (rd_data),   // ?i???????`??
		.rdy_	  (rdy_),	   // ????
		/********** Interrupt  **********/
		.irq_rx	  (irq_rx),	   // ???????????z??
		.irq_tx	  (irq_tx),	   // ???????????z??
		/********** ??????? **********/
		// ????????
		.rx_busy  (rx_busy),   // ?????刅??
		.rx_end	  (rx_end),	   // ???????????
		.rx_data  (rx_data),   // ?????`??
		// ????????
		.tx_busy  (tx_busy),   // ?????刅??
		.tx_end	  (tx_end),	   // ???????????
		.tx_start (tx_start),  // ?????_????
		.tx_data  (tx_data)	   // ?????`??
	);

	/********** UART???????`?? **********/
	uart_tx uart_tx (
		/********** ????a? & ???a? **********/
		.clk	  (clk),	   // ????a?
		.reset	  (reset),	   // ???????a?
		/********** ??????? **********/
		.tx_start (tx_start),  // ?????_????
		.tx_data  (tx_data),   // ?????`??
		.tx_busy  (tx_busy),   // ?????刅??
		.tx_end	  (tx_end),	   // ???????????
		/********** Transmit Signal **********/
		.tx		  (tx)		   // UART???????
	);

	/********** UART???????`?? **********/
	uart_rx uart_rx (
		/********** ????a? & ???a? **********/
		.clk	  (clk),	   // ????a?
		.reset	  (reset),	   // ???????a?
		/********** ??????? **********/
		.rx_busy  (rx_busy),   // ?????刅??
		.rx_end	  (rx_end),	   // ???????????
		.rx_data  (rx_data),   // ?????`??
		/********** Receive Signal **********/
		.rx		  (rx)		   // UART???????
	);

endmodule
