﻿/*
 -- ============================================================================
 -- FILE NAME	: spm.v
 -- DESCRIPTION : spm RAM模块
 -- ----------------------------------------------------------------------------
 -- Revision  Date		  Coding_by	 Comment
 -- 1.0.0	  2011/06/27  suito		 ??????? 
 -- ============================================================================
*/

/********** 通用头文件 **********/
`include "nettype.h"
`include "global_config.h"
`include "stddef.h"

/********** 模块头文件**********/
`include "spm.h"

/********** 模块 **********/
module spm (
	/********** 输入输出参数 **********/
	input  wire				   clk,				// 时钟
	/********** 端口A : IF阶段 **********/
	input  wire [`SpmAddrBus]  if_spm_addr,		// ?????
	input  wire				   if_spm_as_,		// ??????????`??
	input  wire				   if_spm_rw,		// ?i???????
	input  wire [`WordDataBus] if_spm_wr_data,	// ?????z???`??
	output wire [`WordDataBus] if_spm_rd_data,	// ?i???????`??
	/********** 端口B : MEM阶段 **********/
	input  wire [`SpmAddrBus]  mem_spm_addr,	// ?????
	input  wire				   mem_spm_as_,		// ??????????`??
	input  wire				   mem_spm_rw,		// ?i???????
	input  wire [`WordDataBus] mem_spm_wr_data, // ?????z???`??
	output wire [`WordDataBus] mem_spm_rd_data	// ?i???????`??
);

	/********** ?????z???????? **********/
	reg						   wea;			// ??`?? A
	reg						   web;			// ??`?? B

	/********** ?????z????????????? **********/
	always @(*) begin
		/* 端口A */
		if ((if_spm_as_ == `ENABLE_) && (if_spm_rw == `WRITE)) begin   
			wea = `MEM_ENABLE;	// ?????z?????
		end else begin
			wea = `MEM_DISABLE; // ?????z??o??
		end
		/* 端口B */
		if ((mem_spm_as_ == `ENABLE_) && (mem_spm_rw == `WRITE)) begin
			web = `MEM_ENABLE;	// ?????z?????
		end else begin
			web = `MEM_DISABLE; // ?????z??o??
		end
	end

	/********** Xilinx FPGA Block RAM :->altera_dpram **********/
	altera_dpram x_s3e_dpram (
		/********** 端口A : IF????`?? **********/
		.clock_a  (clk),			  // ????a?
		.address_a (if_spm_addr),	  // ?????
		.data_a  (if_spm_wr_data),  // ?????z???`????????A??
		.wren_a   (wea),			  // ?????z???????????`???
		.q_a (if_spm_rd_data),  // ?i???????`??
		/********** 端口B : MEM????`?? **********/
		.clock_b  (clk),			  // ????a?
		.address_b (mem_spm_addr),	  // ?????
		.data_b  (mem_spm_wr_data), // ?????z???`??
		.wren_b   (web),			  // ?????z?????
		.q_b (mem_spm_rd_data)  // ?i???????`??
	);
  
endmodule
